`timescale 1ps/1ps
module Data_Cache(
    input Clk, 
    input Clk_uart,
    input Resetb,
    input DCE_ReadCache,//read write enable signals
    input SB_WriteCache,
    ///////////////////////////////
    //lw from lsq
    input [4:0] Iss_LdStRobTag,
    input [31:0] Iss_LdStAddr, 
    input [5:0] Iss_LdStPhyAddr, 
    ///////////////////////
    input Cdb_Flush,
    input [4:0] Rob_TopPtr,
    input [4:0] Cdb_RobDepth,
    //////////////////////////////////////////
    input [31:0] SB_AddrDmem,
    input [31:0] SB_DataDmem,
    output reg DCE_Opcode,//to ls buffer, for read operation only
    output reg [4:0] DCE_RobTag, 
    output reg [31:0] DCE_Addr,   
    output [31:0] DCE_MemData ,//不能是register
    output reg [5:0] DCE_PhyAddr,//rd physical register number for lw
    //----------------new pin added for CDB-----------
    output DCE_ReadDone,
    //重点：去掉了addr[5:2]=0时直接cache hit的情况，现将延时存入counter再产生done信号，至少一个clock的延时，从而打破loop
    //lsqswaddr[5:2]->read_done->ready-issue->issue addr->lsqswaddr
    output reg DCE_WriteDone,
    output reg DCE_ReadBusy,
    //read busy signal is generated by ls buffer
    output reg DCE_WriteBusy ,
    input Cache_Init, //state signal for initializing data cache
    input Send_DataBack,//state signal for sending data back
    input Uart_DataCache_WE,
    input [5:0] Uart_Cache_InitAddr,//data cache and inst cache can share the same write address for initialization
    input [5:0] Uart_DataCache_RdAddr, 
    input [31:0] Uart_Cache_InitData,
    output [31:0] DataCache_BackData
);
    // parameter File_Name="data_cache_initialization.txt";
    //////////////////////////////////////////////////////////////////////
    //由于设立了SAB，这保证data cache可以同时处理读写操作，但是这里的cache并不是真是的，因此虽然lw,sw的32bit address不同，但是他们【7:2】可能是相同的，
    //测试时应该避免这种情况出现，因为真实cache中，并不只是通过【7:2】address进行写入，这里只是为了简化代码
    //////////////////////////////////////////////////////////////////////
    reg [3:0] LW_Latency_Cnt;//由于访问地址都是提取一个word，因此后两位地址时钟是00，因此将[5:2]4bit用于模拟access latency
    reg [3:0] SW_Latency_Cnt;
    //////////////////////////////////////////////////////////
    ////////////////////////////////////////////////////////
    wire DCE_Flush;
    assign DCE_Flush=(Cdb_Flush&&DCE_RobTag-Rob_TopPtr>Cdb_RobDepth)?1'b1:1'b0;
    //this module is considered as part of tb
    // reg [31:0] Cache_RAM [63:0];
    wire [5:0] wr_addr, rd_addr;
    wire [31:0] din, dout;
    reg write_en;
    /////////////////////////////////
    //clock signals after global mux
    wire Clk2DC_Bram;
    BUFGMUX BUFGMUX_DC (
    .O(Clk2DC_Bram),   // 1-bit output: Clock output
    .I0(Clk), // 1-bit input: Clock input (S=0)
    .I1(Clk_uart), // 1-bit input: Clock input (S=1)
    .S(Cache_Init|Send_DataBack)    // 1-bit input: Clock select
    );
    ///////////////////////////////////
    //memory control signals afer mux
    wire DataCache_WE;
    wire [31:0] DataCache_Din, DataCache_Dout;
    wire [5:0] DataCache_WrAddr, DataCache_RdAddr;

    assign DataCache_WE=Cache_Init?Uart_DataCache_WE:write_en;
    assign DataCache_Din=Cache_Init?Uart_Cache_InitData:SB_DataDmem;
    assign DataCache_WrAddr=Cache_Init?Uart_Cache_InitAddr:SB_AddrDmem[7:2];
    assign DataCache_RdAddr=Send_DataBack?Uart_DataCache_RdAddr:DCE_Addr[7:2];
    //data cache output port assignment 
    assign DCE_MemData=DataCache_Dout;
    assign DataCache_BackData=DataCache_Dout;
    //simple Dual port RAM instantiate
    // dist_mem_gen_1 Cache_RAM (
    // .a(SB_AddrDmem[7:2]),        // input wire [5 : 0] a
    // .d(SB_DataDmem),        // input wire [31 : 0] d
    // .dpra(DCE_Addr[7:2]),  // input wire [5 : 0] dpra
    // .clk(Clk),    // input wire clk
    // .we(write_en),      // input wire we
    // .dpo(DCE_MemData)    // output wire [31 : 0] dpo
    // );
    Uart_Bram Cache_Bram(
        .clk(Clk2DC_Bram),
        .we(DataCache_WE),
        .din(DataCache_Din),//write data in
        .addra(DataCache_WrAddr),//port for write
        .addrb(DataCache_RdAddr),//port for read
        .dout(DataCache_Dout)
    );
    // initial begin
    //     $readmemh(File_Name,Cache_RAM); 
    // end
    //read operation
    ///////////////////////////////////////
    always@(posedge Clk, negedge Resetb)begin
        if(!Resetb)begin
            LW_Latency_Cnt<='bx;
            DCE_RobTag<='bx; 
            DCE_Addr<='bx;
            DCE_PhyAddr<='bx;
            DCE_ReadBusy<=1'b0;
            DCE_Opcode<=1'bx;
        end else begin
            //如果当前时钟发送一个lw,但是被flush掉了，那么这个lw的issue信号根本不会激活，所以当ready cache激活时，不需要考虑cdb flush的影响
            if(!DCE_ReadBusy&&DCE_ReadCache)begin
                DCE_ReadBusy<=!DCE_ReadBusy;
                DCE_RobTag<=Iss_LdStRobTag; 
                DCE_Addr<=Iss_LdStAddr;
                DCE_PhyAddr<=Iss_LdStPhyAddr;
                DCE_Opcode<=DCE_ReadCache;
                if(Iss_LdStAddr[5:2]!=4'b0000)begin
                    LW_Latency_Cnt<=Iss_LdStAddr[5:2];
                end else begin
                    LW_Latency_Cnt<='b1;;//read modified for one clock delay of reading a bram
                end
            end else if(DCE_ReadBusy)begin
                if(DCE_Flush)begin
                    DCE_ReadBusy<=!DCE_ReadBusy;
                end else begin
                    if(LW_Latency_Cnt==4'b0000)begin
                         DCE_ReadBusy<=!DCE_ReadBusy;
                    end else begin
                        LW_Latency_Cnt<=LW_Latency_Cnt-1;
                    end  
                end    
            end
        end
    end
    //重点：原本的计划是用address的最后几bit模拟延时，但是为了仿真无cache miss的情况，是read done是一个纯组合逻辑，但是存在timing loop,
    //为了打破loop，只能将read done改为至少拥有一个clock的延时，但是真时中的cache显然是可以实现cache hit，即无延时读取的，但这里不可以
    //////////////////////////////////////
    //generate read done and read out data
    assign DCE_ReadDone=!DCE_Flush&&DCE_ReadBusy&&LW_Latency_Cnt==4'b0000;  
    ///////////////////////////////////////////////////////////////////////
    //write operation
    always@(posedge Clk, negedge Resetb)begin
        if(!Resetb)begin
            DCE_WriteBusy=1'b0;
            SW_Latency_Cnt<='bx;
        end else begin
            if(SB_WriteCache&&!DCE_WriteBusy)begin
                if(SB_AddrDmem[5:2]!=4'b0000)begin
                    SW_Latency_Cnt<=SB_AddrDmem[5:2]-1;
                    DCE_WriteBusy<=~ DCE_WriteBusy;
                end 
            end
            if(DCE_WriteBusy)begin
                if(SW_Latency_Cnt>0)begin
                    SW_Latency_Cnt<=SW_Latency_Cnt-1;
                end else begin
                    DCE_WriteBusy<=~DCE_WriteBusy;
                    // Cache_RAM[SB_AddrDmem[7:2]]<=SB_DataDmem;
                end
            end
        end
    end
    //////////////////////////////////////////////////
    always@(*)begin
        DCE_WriteDone=1'b0;
        write_en=1'b0;
        if(SB_WriteCache&&!DCE_WriteBusy&&SB_AddrDmem[5:2]==4'b0000)begin
            DCE_WriteDone=1'b1;
            write_en=1'b1;
        end else if(DCE_WriteBusy&&SW_Latency_Cnt==4'b0000)begin
            DCE_WriteDone=1'b1;
            write_en=1'b1;
        end
    end
    
endmodule